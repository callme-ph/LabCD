entity Or3In is
	port(
		entry1, entry2, entry3: in bit;
		or_out: out bit
	);
end Or3In;

architecture behav of Or3In is

begin
	or_out <= entry1 or entry2 or entry3;
	
end architecture behav;