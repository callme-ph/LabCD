library verilog;
use verilog.vl_types.all;
entity Lab02_vlg_check_tst is
    port(
        s1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab02_vlg_check_tst;
