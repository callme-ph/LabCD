library verilog;
use verilog.vl_types.all;
entity Lab02 is
    port(
        s1              : out    vl_logic;
        c               : in     vl_logic;
        b               : in     vl_logic;
        a               : in     vl_logic
    );
end Lab02;
