library verilog;
use verilog.vl_types.all;
entity Lab02_vlg_vec_tst is
end Lab02_vlg_vec_tst;
